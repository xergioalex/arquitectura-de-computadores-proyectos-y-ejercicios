library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Logica is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           C : out  STD_LOGIC);
end Logica;

architecture Behavioral of Logica is

begin


end Behavioral;

