library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Compuerta is
end Compuerta;

architecture Behavioral of Compuerta is

begin


end Behavioral;

