`timescale 1ns / 1ps

module algoc(
	 input a,
	 input b,
	 output so
	 );
	 assing so = a ^ b;

endmodule
